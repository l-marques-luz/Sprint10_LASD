module clock1s(
input clock,
output reg clocknovo
);
reg [25:0] contador;
always @(posedge clock)
begin
	if (contador == 25000000/10) 
	begin
		clocknovo = ~clocknovo;
		contador = 0;
	end
	else
	contador = contador + 1;
end
endmodule